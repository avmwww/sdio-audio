// TDM front end

module tdm_fe(
	input  wire        iclk,
	input  wire        irst,
	input  wire [31:0] idata,	// Input data
	input  wire        idata_en,	// Input data enable
	input  wire        iout_data_dis,// disable output data
	output wire [31:0] odata,	// Output data
	output wire        odata_en,	// Output data enable
);

endmodule
