// Clock generation module

module clk_rst_gen(
	output wire oclk, // generated lock
	output wire orst  // generated reset
);


endmodule
