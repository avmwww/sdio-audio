// Verification module


module verif(
	input  wire imclk,  // Master clock input
	input  wire ifs,    // Frame sync
	input  wire isclk,  // Serial clock
	input  wire idin,   // Serial data input
	output wire odout   // Serial data output
);

endmodule
