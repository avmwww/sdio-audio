// TDM serializer

module tdm_sh(
	input  wire        iclk,
	input  wire        irst,
	input  wire [31:0] idata,
	output wire        odata_en,
	output wire        odout
);

endmodule

