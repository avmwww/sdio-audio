// TDM serializer

module tdm_sh(
);

endmodule
