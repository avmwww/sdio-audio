// TDM back end

module tdm_be(
	input  wire        iclk,
	input  wire        irst,
	input  wire [31:0] idin,	// Input data
	output wire        odin_en,	// Input data enable
	input  wire        idout_en,	// Output data enable
	output wire [31:0] odout,	// Output data
);

endmodule
